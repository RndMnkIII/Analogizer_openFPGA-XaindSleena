//xain_top.sv
